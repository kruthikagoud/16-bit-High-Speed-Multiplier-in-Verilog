`timescale 1 ns / 1 ns
module mul16(a,b,o);
input [15:0]a,b;
output [31:0]o;
wire [31:0]o1,o2,o3,o4,o5,o6,o7,o8,o9,o10,o11,o12,o13,o14,o15,o16;
assign o1=b[0]?({16'b0000000000000000,a[15:0]}):32'b00000000000000000000000000000000;
assign o2=b[1]?({15'b000000000000000,a[15:0],1'b0}):32'b00000000000000000000000000000000;
assign o3=b[2]?({14'b00000000000000,a[15:0],2'b00}):32'b00000000000000000000000000000000;
assign o4=b[3]?({13'b0000000000000,a[15:0],3'b000}):32'b00000000000000000000000000000000;
assign o5=b[4]?({12'b000000000000,a[15:0],4'b0000}):32'b00000000000000000000000000000000;
assign o6=b[5]?({11'b00000000000,a[15:0],5'b00000}):32'b00000000000000000000000000000000;
assign o7=b[6]?({10'b0000000000,a[15:0],6'b000000}):32'b00000000000000000000000000000000;
assign o8=b[7]?({9'b000000000,a[15:0],7'b0000000}):32'b00000000000000000000000000000000;
assign o9=b[8]?({8'b00000000,a[15:0],8'b00000000}):32'b00000000000000000000000000000000;
assign o10=b[9]?({7'b0000000,a[15:0],9'b000000000}):32'b00000000000000000000000000000000;
assign o11=b[10]?({6'b000000,a[15:0],10'b0000000000}):32'b00000000000000000000000000000000;
assign o12=b[11]?({5'b00000,a[15:0],11'b00000000000}):32'b00000000000000000000000000000000;
assign o13=b[12]?({4'b0000,a[15:0],12'b000000000000}):32'b00000000000000000000000000000000;
assign o14=b[13]?({3'b000,a[15:0],13'b0000000000000}):32'b00000000000000000000000000000000;
assign o15=b[14]?({2'b00,a[15:0],14'b00000000000000}):32'b00000000000000000000000000000000;
assign o16=b[15]?({1'b0,a[15:0],15'b000000000000000}):32'b00000000000000000000000000000000;
assign o = o1+o2+o3+o4+o5+o6+o7+o8+o9+o10+o11+o12+o13+o14+o15+o16;
endmodule



module mul16_tb;
reg [15:0]a,b;
wire [31:0]o;
mul16 a1(a,b,o);
initial
repeat(10)
begin
a=$random;
b=$random;
#100;
end
endmodule
